


#        ScrollAnywhere
app_name=ScrollAnywhere
#        Drag scrollbar with your middle mouse button anywhere on the page. Supports also "grab and drag" style and Momentum.
app_desc=Dra rullningslisten med din mittmusknapp var som helst på sidan. Stöder även "ta och dra" och rörelsemängd.

#                       Default value: $1, min: $2, max: $3
field_int_default_value=Standardvärde: $1, min: $2, max: $3
#                 Reset to default: $1
field_set_default=Återställ till standard: $1


#                 Thunderbird Add-ons page
thunderbird_store=
#             Firefox Add-ons page
firefox_store=Firefox tilläggssida
#            Chrome Web Store page
chrome_store=Chrome Web Store-sidan
#           Disable on $1
win_disable=Inaktiverad på $1
#                                Disable horizontal scrolling on $1
win_horizontal_scrolling_disable=
#             Visit homepage
op_visit_home=Besök hemsidan
#             Help this project
op_support_me=Hjälp det här projektet


#       Options - $1
o_title=Alternativ - $1
#             General
o_tab_general=Allmänt
#              Momentum
o_tab_momentum=Rörelsemängd
#            Cursor
o_tab_cursor=Markör
#              Axis locking
o_axis_locking=
#                 Performance
o_tab_performance=Prestanda
#                 Disabled on
o_tab_disabled_on=Inaktiverad på
#              Advanced
o_tab_advanced=Avancerat
#                Scrollbars
o_tab_scrollbars=
#            Backup
o_tab_backup=Säkerhetskopia
#           About
o_tab_about=Om

#                  When scrolling a box that is scrollable in one axis but parent box is scrollable in other axis, lock scrolling to one axis using:
o_axis_lock_helper=
#             Smart lock - temporal lock using momentum
o_axis_lock_0=
#             Strict lock - instant direction lock
o_axis_lock_1=
#             No lock - free scrolling in both axis
o_axis_lock_2=
#                       Smart lock stack size
o_trend_momentum_window=
#                              Larger value will require more scrolling in opposite axis to change the scrolling axis.
o_trend_momentum_window_helper=

#                        Addon is disabled! Click here to enable.
o_addon_disabled_warning=

#                       no change - best performance
o_cursor_change_default=ingen ändring - bästa prestanda
#               Scroll button:
o_scroll_button=Rullningsknapp:
#                 Scroll style  / direction / speed:
o_direction_speed=Rullningsstil / riktning / hastighet:
#            Multiplier
o_multiplier=Multiplikator
#             times scroll speed
o_times_speed=gånger rullhastighet

#               Maximum scroll speed (0 - disabled):
o_maximum_speed=Maximal rullhastighet (0 - inaktiverad):
#            ratio (page length / window size)
o_ratio_unit=förhållande (sidlängd / fönsterstorlek)

#               Emulate Scrollbar
o_scroll_type_0=Emulera rullningslist
#               Grab and Drag - like on a smartphone
o_scroll_type_1=Ta och dra - som på en smartmobil
#               Dynamic Speed (experimental)
o_scroll_type_2=Dynamisk hastighet (experimentell)
#                     It's like dragging a scrollbar
o_scroll_type_title_0=Det är som att dra en rullningslist
#                     It's like dragging a page with your finger on a phone screen
o_scroll_type_title_1=Det är som att dra en sida med ditt finger på en telefonskärm
#                     Dynamic Speed makes scroll speed slower when page is longer
o_scroll_type_title_2=Dynamisk hastighet gör rullhastigheten långsammare när sidan är längre

#             Disable / Enable scrolling when key is down:
o_disable_key=Inaktivera / Aktivera rullning när tangent hålls nertryckt:
#                   Momentum:
o_momentum_category=Rörelsemängd:

#                  Momentum formula:
o_momentum_formula=Rörelseformel:
#                         Uniformly decelerated movement
o_momentum_formula_type_0=Likformig hastighetsmindskningsrörelse
#                               Page scroll will be uniformly slowed down until it stops
o_momentum_formula_type_title_0=Sidrullning kommer att med jämn hastighet sänkas tills tills den stannar helt
#                         Exponentially decelerated movement
o_momentum_formula_type_1=Exponentiellt decelererad rörelse
#                               Page scroll will rapidly (exponentially) slow down
o_momentum_formula_type_title_1=Sidrullning kommer snabbt (exponentiellt) att sänkas
#                         Infinite movement ∞
o_momentum_formula_type_2=Oändlig rörelse ∞
#                               Scrolling will never stop
o_momentum_formula_type_title_2=Rullningen kommer aldrig stanna

#                    Maximum speed (0 - disabled):
o_momentum_max_speed=Max hastighet (0 - inaktiverad):

#             Page weight:
o_page_weight=Sidvikt:
#       grams :)
o_grams=gram :)
#                  Additional speed:
o_additional_speed=Ytterliggare hastighet:
#               pixels per second
o_pixels_second=pixlar per sekund
#                     Additional duration:
o_additional_duration=Ytterligare varaktighet:
#              milliseconds
o_milliseconds=millisekunder
#                   Advanced momentum setup (for experts only!):
o_advanced_momentum=Avancerad rörelsemängdinställning (endast för experter!):
#                         Changing these values can break your momentum!
o_advanced_momentum_title=Ändras dessa värden kan rörelsemängden sluta fungera!
#                   Compute from last:
o_compute_from_last=Beräkna från sista:
#                      Mouse stop detection:
o_mouse_stop_detection=Musstoppsdetektering:
#                Tracking speed:
o_tracking_speed=Spårhastighet:
#              Reset values
o_reset_values=Återställ värden
#                  Cursor used when scrolling:
o_cursor_scrolling=Markör som används när du rullar:
#             Performance:
o_performance=Prestanda:
#                   Prevent big jumps
o_prevent_big_jumps=
#                          If you are using tool that can teleport your cursor across the screen (when you reach an edge), enable this option to allow continuous (infinite) scrolling.
o_prevent_big_jumps_helper=
#          Advanced:
o_advanced=Avancerat:
#                    Mouse movement detection threshold:
o_movement_detection=Detektionsgränsen för musrörelse:
#                            How many pixels has to mouse move to block link. Sometimes when pressing scroll button you move mouse slightly but you don't want the link to be disabled because of that.
o_helper_text_move_detection=Hur många pixlar måste musen flytta sig för att blockera länkar. Ibland när du trycker på rullningsknappen flyttar du musen litegrann, men du vill inte att länken ska inaktiveras på grund av det.
#                    Context menu block:
o_context_menu_block=
#                            Unblock context menu delay
o_context_menu_unblock_delay=
#                                   If you see context menu after scrolling with Right mouse button, increase this value
o_context_menu_unblock_delay_helper=

#       times
o_times=gånger
#        pixels
o_pixels=pixlar
#       items
o_items=

#                                       Disable horizontal scrolling on domains:
o_disabled_horizontal_scrolling_domains=
#                     Disabled on domains:
o_is_disabled_domains=Inaktiverad på domäner:
#                 Disabled on pages / sub-pages:
o_is_disabled_url=Inaktiverad på sidor / undersidor:
#                      You can use star symbol (*) to define a URL part, for example: "google.com/maps*"
o_is_disabled_url_help=Du kan använda en asterisk (*) för att definiera en del av en webbadress, till exempel: "google.se/maps*"
#             Disable add-on
o_is_disabled=Inaktivera tillägg
#                      Middle button
o_scroll_button_middle=Mittknapp
#                     Right button
o_scroll_button_right=Högerknapp
#                                Linux / Mac users - you will be prompted for new permission "Read and modify browser setting" - this is required to suppress context menu being shown before scrolling!
o_scroll_button_right_linux_note=Linux- / Mac-användare - du kommer att bli tillfrågan om en ny behörighet "Läs och ändra webbläsarinställningar" - detta krävs för att förhindra att innehållsmenyn visas före du rullar!
#                                       Linux / Mac users - your context menu will be blocked! To open context menu hold "Shift" key or triple-click right button.
o_scroll_button_right_linux_chrome_note=Linux- / Mac-användare - din innehållsmeny kommer att blockeras! För att öppna innehållsmenyn håller du knappen "Skift" nertryckt eller trippelklickar på högerknappen.
#                    Left button (experimental)
o_scroll_button_left=Vänsterknapp (experimentell)
#                 Scroll on links
o_scroll_on_links=Rulla på länkar
#                       When enabled, you won't be able to drag and drop links (only by using 'Disable' key)
o_scroll_on_links_title=När detta är aktiverat kommer du inte att kunna dra och släppa länkar (endast om "Inaktivera"-tangenten används)
#                Scroll on text
o_scroll_on_text=
#                      Emulates phone scrolling / editing - you need to click on text in order to switch to "editing mode". Clicking outside of text enables scrolling again.
o_scroll_on_text_title=
#                    Scroll on textarea
o_scroll_on_textarea=
#                          Textarea is a block of text, usually resizable. For example on "Disabled on" tab you can see textarea.
o_scroll_on_textarea_title=
#                         Scroll on editable html
o_scroll_on_editable_html=
#                               For example email body in Gmail is editable html.
o_scroll_on_editable_html_title=

#                          on text will enable selecting / editing text.
o_scroll_on_text_edit_with=
#                                Click on text will enable "Edit mode". Click outside text to enable "Scroll mode".
o_scroll_on_text_edit_with_title=
#                            Single click
o_scroll_on_text_edit_with_0=
#                            Double click
o_scroll_on_text_edit_with_1=

#                  Scrollbars look
o_scrollbars_width=
#                    Normal (no change)
o_scrollbars_width_0=
#                    Thin
o_scrollbars_width_1=
#                    Hidden
o_scrollbars_width_2=

#                  Scrollbar slider color:
o_scrollbars_color=
#                       Scrollbar background color:
o_scrollbars_background=

#         Reverse scroll direction
o_reverse=Omvänd rullningsriktning
#             Alt
o_disable_alt=Alt
#               Shift
o_disable_shift=Skift
#              Ctrl
o_disable_ctrl=Ctrl
#                Disable when key is down:
o_disable_type_0=Inaktivera när tangent hålls nertryckt:
#                Enable when key is down:
o_disable_type_1=Aktivera när tangent hålls nertryckt:
#          disabled
o_disabled=inaktiverad
#         enabled
o_enabled=aktiverad
#          enable momentum - you can "throw" the page (like on phone)
o_momentum=aktivera momentum - du kan "kasta" sidan (som på en pektelefon)
#             Don't lock iframes and don't change cursor when scrolling
o_no_css_edit=Lås inte iframes och ändra inte markören när du rullar
#                    Don't block default button action
o_no_prevent_default=Blockera inte standardknappsåtgärd
#                Links blocking:
o_auto_link_lock=Link blockering:
#               Don't block mouse click on link after movement
o_no_link_block=Blockera inte musklick på länken efter rörelse
#                               When you start scrolling on a link and then you finish scrolling on the same link, browser will open the link. This is usually not desired behaviour so by default it's blocked.
o_helper_text_middle_link_click=När du börjar rulla på en länk och du sedan slutar rulla på samma länk, då öppnar webbläsaren länken. Detta är vanligtvis inte ett önskat beteende så detta är blockerat som standard.

#                   This controls how 'heavy' the page is. Heavier pages has longer momentum.
o_page_weight_title=Detta kontrollerar hur "tung" sidan är. Tyngre sidor har längre rörelsemängd.
#                        You can accelerate momentum stating speed.
o_additional_speed_title=Du kan accelerera hastigheten på rörelsemängden.
#                           Additional time for each momentum.
o_additional_duration_title=Ytterliggare tid för varje rörelsemängd.
#                         Momentum initial speed is determined by the speed of scrolling right before releasing the Scroll button.
o_compute_from_last_title=Rörelsemängdens initialhastighet avgörs av rullhastigheten precis innan du släpper rullknappen.
#                            How much time has to mouse stay still - before releasing the Scroll button - to NOT activate Momentum.
o_mouse_stop_detection_title=Hur mycket tid måste musen stå still - innan du släpper rullningsknappen - för att INTE aktivera rörelsemängd.
#                      Interval for measuring current scroll speed.
o_tracking_speed_title=Intervall för mätning av aktuell rullhastighet.
#                Scrolling area:
o_scrolling_area=
#                    Scrolling area (0 - disabled):
o_outside_area_width=
#                           Moving your cursor outside of scrolling area will revert scrolling position. Same behavior can be seen when dragging a scrollbar.
o_outside_area_width_helper=

#                          Warning - Left button support is using deprecated Firefox API that could be removed in future versions of Firefox.
o_scroll_button_left_title=Varning - Vänster knappstöd använder vanligt Firefox-API som kan tas bort i framtida versioner av Firefox.
#                        Prevent text selection when scrolling with left button
o_prevent_text_selection=Förhindra att text markeras när du rullar med vänster knapp
#                                    On some devices, scrolling with left mouse button will also select text on the page.
o_helper_text_prevent_text_selection=På vissa enheter kommer texten att markeras när du använder vänster musknapp att rulla med.

#                              Don't block context menu when trying to scroll not-scrollable page
o_disable_context_menu_on_move=Blockera inte innehållsmenyn när du försöker rulla på en icke-rullbar sida


#                Backup / Restore settings:
o_backup_restore=Säkerhetskopiera / Återställ inställningar:
#                 Export settings to a file
o_export_settings=Exportera inställningar till en fil
#                      Import settings from $1 file...
import_settings_button=Importera inställningar från filen $1 ...
#               Import finished!
import_finished=Importerad!
#             working...
label_working=arbetar...


#               Test your scrolling settings here
test_page_title=Testa dina rullningsinställningar här


#            Options
menu_options=Alternativ
#                Visit homepage
menu_visit_title=Besök hemsida
#           Disabled by your web-browser
not_working=Inaktiverad av din webbläsare
#                Disabled on this domain
disabled_by_user=
#                 Your browser will block ScrollAnywhere on these type of pages:
not_working_title=Din webbläsare blockerar ScrollAnywhere på dessa typer av sidor:
#                To enable ScrollAnywhere on "mozilla.org" pages, see this YouTube tutorial
not_working_body=För att aktivera ScrollAnywhere på sidor som "mozilla.org", titta på denna handledning på YouTube

#           Close
label_close=Stäng


#             Switch add-on OFF / ON
switch_on_off=Växla tillägget AV / PÅ

#                                If you experience noticeable delay between pressing scroll button and starting scrolling, try to enable this option. However you will not be able to scroll over "iframes" such as some old embedded videos or some ads.
o_helper_text_performance_iframe=Om du upplever märkbar fördröjning mellan att trycka på rullningsknappen och starta rullningen, försök aktivera det här alternativet. Du kommer dock inte att kunna rulla över "iframes" som en del gamla inbäddade videor eller annonser.
#                                This will also disable option to change cursor while scrolling.
o_helper_text_performance_cursor=Detta kommer också att inaktivera alternativet att byta markör medan du bläddrar.
#                            Useful in Linux to enable Paste with middle button.
o_helper_text_default_action=Användbar i Linux för att aktivera "Klistra in" med mittknappen.

#             Hello :)
o_about_hello=Hej :)
#             My name is Juraj Mäsiar and I'm the author of ScrollAnywhere.
o_about_intro=Jag heter Juraj Mäsiar och jag är skaparen av ScrollAnywhere.
#               If you like it, please rate it here:
o_about_like_it=Om du gillar det, betygsätt gärna det här:
#                  If you don't like it, please let me know why to my e-mail. I'm implementing most of the feature-requests I receive.
o_about_dislike_it=Om du inte gillar det, vill jag gärna att du skickar ett e-postmeddelande och talar om varför. Jag genomför de flesta av de funktionsförfrågningar jag får.

#                  Please consider supporting my work by
o_about_support_by=Stöd gärna mitt arbete genom
#                           donation (PayPal)
o_about_support_by_donation=donation (PayPal)
#                         becoming my Patron
o_about_support_by_patron=blir min Patron

#              Thank you!
o_about_thanks=Tack!
#            home:
o_about_home=hem:
#               Contact:
o_about_contact=Kontakta:
#              Report issues:
o_about_issues=
#                     I can reply only in English / Slovak
o_about_support_reply=Jag kan bara svara på Engelska / Slovakiska
#                    Social media:
o_about_social_media=Sociala medier:
#            Save changes and close
o_save_close=Spara ändringar och stäng
#       saved!
o_saved=sparad!


#                 Coming soon
label_coming_soon=Kommer snart
#                  Save changes
label_save_changes=Spara ändringar
